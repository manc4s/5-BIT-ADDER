`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01/25/2025 07:55:04 PM
// Design Name: 
// Module Name: 5bit_addition
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module 5bit_addition(
    input a0,
    input a1,
    input a2,
    input a3,
    input a4,
    input b0,
    input b1,
    input b2,
    input b3,
    input b4,
    output s0,
    output s1,
    output s2,
    output s3,
    output s4,
    input cin,
    output cout
    );
endmodule
